// cTypes = List(3, 4, 3, 3, 4, 4)
module BoothCodeUnit(
  input  [64:0] io_A,
  input  [2:0]  io_code,
  output [65:0] io_boothCodeOutput_product,
  output [1:0]  io_boothCodeOutput_h,
  output        io_boothCodeOutput_sn
);
  wire  A_sign = io_A[64]; // @[BoothCode.scala 23:17]
  wire [65:0] _io_boothCodeOutput_product_T = {A_sign,io_A}; // @[Cat.scala 31:58]
  wire  _io_boothCodeOutput_sn_T = ~A_sign; // @[BoothCode.scala 31:30]
  wire [65:0] _io_boothCodeOutput_product_T_2 = {io_A,1'h0}; // @[Cat.scala 31:58]
  wire [64:0] _io_boothCodeOutput_product_T_3 = ~io_A; // @[BoothCode.scala 42:39]
  wire [65:0] _io_boothCodeOutput_product_T_4 = {_io_boothCodeOutput_product_T_3,1'h1}; // @[Cat.scala 31:58]
  wire [65:0] _io_boothCodeOutput_product_T_7 = {_io_boothCodeOutput_sn_T,_io_boothCodeOutput_product_T_3}; // @[Cat.scala 31:58]
  wire  _T_6 = io_code == 3'h6; // @[BoothCode.scala 49:22]
  wire [65:0] _GEN_3 = io_code == 3'h6 ? _io_boothCodeOutput_product_T_7 : 66'h0; // @[BoothCode.scala 49:36 50:32]
  wire  _GEN_4 = io_code == 3'h6 ? A_sign : 1'h1; // @[BoothCode.scala 49:36 51:27]
  wire [65:0] _GEN_6 = io_code == 3'h5 ? _io_boothCodeOutput_product_T_7 : _GEN_3; // @[BoothCode.scala 45:36 46:32]
  wire  _GEN_7 = io_code == 3'h5 ? A_sign : _GEN_4; // @[BoothCode.scala 45:36 47:27]
  wire  _GEN_8 = io_code == 3'h5 | _T_6; // @[BoothCode.scala 45:36 48:26]
  wire [65:0] _GEN_9 = io_code == 3'h4 ? _io_boothCodeOutput_product_T_4 : _GEN_6; // @[BoothCode.scala 41:36 42:32]
  wire  _GEN_10 = io_code == 3'h4 ? A_sign : _GEN_7; // @[BoothCode.scala 41:36 43:27]
  wire  _GEN_11 = io_code == 3'h4 | _GEN_8; // @[BoothCode.scala 41:36 44:26]
  wire [65:0] _GEN_12 = io_code == 3'h3 ? _io_boothCodeOutput_product_T_2 : _GEN_9; // @[BoothCode.scala 37:36 38:32]
  wire  _GEN_13 = io_code == 3'h3 ? _io_boothCodeOutput_sn_T : _GEN_10; // @[BoothCode.scala 37:36 39:27]
  wire  _GEN_14 = io_code == 3'h3 ? 1'h0 : _GEN_11; // @[BoothCode.scala 37:36 40:26]
  wire [65:0] _GEN_15 = io_code == 3'h2 ? _io_boothCodeOutput_product_T : _GEN_12; // @[BoothCode.scala 33:36 34:32]
  wire  _GEN_16 = io_code == 3'h2 ? _io_boothCodeOutput_sn_T : _GEN_13; // @[BoothCode.scala 33:36 35:27]
  wire  _GEN_17 = io_code == 3'h2 ? 1'h0 : _GEN_14; // @[BoothCode.scala 33:36 36:26]
  wire [65:0] _GEN_18 = io_code == 3'h1 ? _io_boothCodeOutput_product_T : _GEN_15; // @[BoothCode.scala 29:36 30:32]
  wire  _GEN_19 = io_code == 3'h1 ? ~A_sign : _GEN_16; // @[BoothCode.scala 29:36 31:27]
  wire  _GEN_20 = io_code == 3'h1 ? 1'h0 : _GEN_17; // @[BoothCode.scala 29:36 32:26]
  wire  _GEN_23 = io_code == 3'h0 ? 1'h0 : _GEN_20; // @[BoothCode.scala 25:30 28:26]
  assign io_boothCodeOutput_product = io_code == 3'h0 ? 66'h0 : _GEN_18; // @[BoothCode.scala 25:30 26:32]
  assign io_boothCodeOutput_h = {{1'd0}, _GEN_23};
  assign io_boothCodeOutput_sn = io_code == 3'h0 | _GEN_19; // @[BoothCode.scala 25:30 27:27]
endmodule
module Compressor32(
  input  [72:0] io_in_0,
  input  [72:0] io_in_1,
  input  [72:0] io_in_2,
  output [72:0] io_s,
  output [72:0] io_ca
);
  wire [72:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [72:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [72:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [72:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [72:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor32_10(
  input  [68:0] io_in_0,
  input  [68:0] io_in_1,
  input  [68:0] io_in_2,
  output [68:0] io_s,
  output [68:0] io_ca
);
  wire [68:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [68:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [68:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [68:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [68:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor42(
  input  [74:0] io_p_0,
  input  [74:0] io_p_1,
  input  [74:0] io_p_2,
  input  [74:0] io_p_3,
  output [74:0] io_s,
  output [74:0] io_ca
);
  wire [74:0] xor0 = io_p_0 ^ io_p_1; // @[Compressor42.scala 19:19]
  wire [74:0] _cout_T = xor0 & io_p_2; // @[Compressor42.scala 23:16]
  wire [74:0] _cout_T_1 = ~xor0; // @[Compressor42.scala 23:30]
  wire [74:0] _cout_T_2 = _cout_T_1 & io_p_0; // @[Compressor42.scala 23:44]
  wire [74:0] cout = _cout_T | _cout_T_2; // @[Compressor42.scala 23:26]
  wire [74:0] cin = {cout[73:0],1'h0}; // @[Cat.scala 31:58]
  wire [74:0] xor1 = io_p_2 ^ io_p_3; // @[Compressor42.scala 20:19]
  wire [74:0] xor2 = xor1 ^ xor0; // @[Compressor42.scala 21:16]
  wire [74:0] _io_ca_T = xor2 & cin; // @[Compressor42.scala 25:17]
  wire [74:0] _io_ca_T_1 = ~xor2; // @[Compressor42.scala 25:27]
  wire [74:0] _io_ca_T_2 = _io_ca_T_1 & io_p_3; // @[Compressor42.scala 25:41]
  assign io_s = xor2 ^ cin; // @[Compressor42.scala 24:16]
  assign io_ca = _io_ca_T | _io_ca_T_2; // @[Compressor42.scala 25:23]
endmodule
module Compressor42_1(
  input  [79:0] io_p_0,
  input  [79:0] io_p_1,
  input  [79:0] io_p_2,
  input  [79:0] io_p_3,
  output [79:0] io_s,
  output [79:0] io_ca
);
  wire [79:0] xor0 = io_p_0 ^ io_p_1; // @[Compressor42.scala 19:19]
  wire [79:0] _cout_T = xor0 & io_p_2; // @[Compressor42.scala 23:16]
  wire [79:0] _cout_T_1 = ~xor0; // @[Compressor42.scala 23:30]
  wire [79:0] _cout_T_2 = _cout_T_1 & io_p_0; // @[Compressor42.scala 23:44]
  wire [79:0] cout = _cout_T | _cout_T_2; // @[Compressor42.scala 23:26]
  wire [79:0] cin = {cout[78:0],1'h0}; // @[Cat.scala 31:58]
  wire [79:0] xor1 = io_p_2 ^ io_p_3; // @[Compressor42.scala 20:19]
  wire [79:0] xor2 = xor1 ^ xor0; // @[Compressor42.scala 21:16]
  wire [79:0] _io_ca_T = xor2 & cin; // @[Compressor42.scala 25:17]
  wire [79:0] _io_ca_T_1 = ~xor2; // @[Compressor42.scala 25:27]
  wire [79:0] _io_ca_T_2 = _io_ca_T_1 & io_p_3; // @[Compressor42.scala 25:41]
  assign io_s = xor2 ^ cin; // @[Compressor42.scala 24:16]
  assign io_ca = _io_ca_T | _io_ca_T_2; // @[Compressor42.scala 25:23]
endmodule
module Compressor42_5(
  input  [75:0] io_p_0,
  input  [75:0] io_p_1,
  input  [75:0] io_p_2,
  input  [75:0] io_p_3,
  output [75:0] io_s,
  output [75:0] io_ca
);
  wire [75:0] xor0 = io_p_0 ^ io_p_1; // @[Compressor42.scala 19:19]
  wire [75:0] _cout_T = xor0 & io_p_2; // @[Compressor42.scala 23:16]
  wire [75:0] _cout_T_1 = ~xor0; // @[Compressor42.scala 23:30]
  wire [75:0] _cout_T_2 = _cout_T_1 & io_p_0; // @[Compressor42.scala 23:44]
  wire [75:0] cout = _cout_T | _cout_T_2; // @[Compressor42.scala 23:26]
  wire [75:0] cin = {cout[74:0],1'h0}; // @[Cat.scala 31:58]
  wire [75:0] xor1 = io_p_2 ^ io_p_3; // @[Compressor42.scala 20:19]
  wire [75:0] xor2 = xor1 ^ xor0; // @[Compressor42.scala 21:16]
  wire [75:0] _io_ca_T = xor2 & cin; // @[Compressor42.scala 25:17]
  wire [75:0] _io_ca_T_1 = ~xor2; // @[Compressor42.scala 25:27]
  wire [75:0] _io_ca_T_2 = _io_ca_T_1 & io_p_3; // @[Compressor42.scala 25:41]
  assign io_s = xor2 ^ cin; // @[Compressor42.scala 24:16]
  assign io_ca = _io_ca_T | _io_ca_T_2; // @[Compressor42.scala 25:23]
endmodule
module Compressor32_11(
  input  [86:0] io_in_0,
  input  [86:0] io_in_1,
  input  [86:0] io_in_2,
  output [86:0] io_s,
  output [86:0] io_ca
);
  wire [86:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [86:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [86:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [86:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [86:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor32_12(
  input  [91:0] io_in_0,
  input  [91:0] io_in_1,
  input  [91:0] io_in_2,
  output [91:0] io_s,
  output [91:0] io_ca
);
  wire [91:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [91:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [91:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [91:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [91:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor32_14(
  input  [87:0] io_in_0,
  input  [87:0] io_in_1,
  input  [87:0] io_in_2,
  output [87:0] io_s,
  output [87:0] io_ca
);
  wire [87:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [87:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [87:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [87:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [87:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor32_15(
  input  [114:0] io_in_0,
  input  [114:0] io_in_1,
  input  [114:0] io_in_2,
  output [114:0] io_s,
  output [114:0] io_ca
);
  wire [114:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [114:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [114:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [114:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [114:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor32_16(
  input  [100:0] io_in_0,
  input  [100:0] io_in_1,
  input  [100:0] io_in_2,
  output [100:0] io_s,
  output [100:0] io_ca
);
  wire [100:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [100:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [100:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [100:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [100:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Compressor42_6(
  input  [125:0] io_p_0,
  input  [125:0] io_p_1,
  input  [125:0] io_p_2,
  input  [125:0] io_p_3,
  output [125:0] io_s,
  output [125:0] io_ca
);
  wire [125:0] xor0 = io_p_0 ^ io_p_1; // @[Compressor42.scala 19:19]
  wire [125:0] _cout_T = xor0 & io_p_2; // @[Compressor42.scala 23:16]
  wire [125:0] _cout_T_1 = ~xor0; // @[Compressor42.scala 23:30]
  wire [125:0] _cout_T_2 = _cout_T_1 & io_p_0; // @[Compressor42.scala 23:44]
  wire [125:0] cout = _cout_T | _cout_T_2; // @[Compressor42.scala 23:26]
  wire [125:0] cin = {cout[124:0],1'h0}; // @[Cat.scala 31:58]
  wire [125:0] xor1 = io_p_2 ^ io_p_3; // @[Compressor42.scala 20:19]
  wire [125:0] xor2 = xor1 ^ xor0; // @[Compressor42.scala 21:16]
  wire [125:0] _io_ca_T = xor2 & cin; // @[Compressor42.scala 25:17]
  wire [125:0] _io_ca_T_1 = ~xor2; // @[Compressor42.scala 25:27]
  wire [125:0] _io_ca_T_2 = _io_ca_T_1 & io_p_3; // @[Compressor42.scala 25:41]
  assign io_s = xor2 ^ cin; // @[Compressor42.scala 24:16]
  assign io_ca = _io_ca_T | _io_ca_T_2; // @[Compressor42.scala 25:23]
endmodule
module Compressor42_7(
  input  [132:0] io_p_0,
  input  [132:0] io_p_1,
  input  [132:0] io_p_2,
  input  [132:0] io_p_3,
  output [132:0] io_s,
  output [132:0] io_ca
);
  wire [132:0] xor0 = io_p_0 ^ io_p_1; // @[Compressor42.scala 19:19]
  wire [132:0] _cout_T = xor0 & io_p_2; // @[Compressor42.scala 23:16]
  wire [132:0] _cout_T_1 = ~xor0; // @[Compressor42.scala 23:30]
  wire [132:0] _cout_T_2 = _cout_T_1 & io_p_0; // @[Compressor42.scala 23:44]
  wire [132:0] cout = _cout_T | _cout_T_2; // @[Compressor42.scala 23:26]
  wire [132:0] cin = {cout[131:0],1'h0}; // @[Cat.scala 31:58]
  wire [132:0] xor1 = io_p_2 ^ io_p_3; // @[Compressor42.scala 20:19]
  wire [132:0] xor2 = xor1 ^ xor0; // @[Compressor42.scala 21:16]
  wire [132:0] _io_ca_T = xor2 & cin; // @[Compressor42.scala 25:17]
  wire [132:0] _io_ca_T_1 = ~xor2; // @[Compressor42.scala 25:27]
  wire [132:0] _io_ca_T_2 = _io_ca_T_1 & io_p_3; // @[Compressor42.scala 25:41]
  assign io_s = xor2 ^ cin; // @[Compressor42.scala 24:16]
  assign io_ca = _io_ca_T | _io_ca_T_2; // @[Compressor42.scala 25:23]
endmodule
module Compressor32_17(
  input  [64:0] io_in_0,
  input  [64:0] io_in_1,
  input  [64:0] io_in_2,
  output [64:0] io_s,
  output [64:0] io_ca
);
  wire [64:0] _io_s_T = io_in_0 ^ io_in_1; // @[Compressor32.scala 21:13]
  wire [64:0] _io_ca_T = io_in_0 & io_in_1; // @[Compressor32.scala 22:15]
  wire [64:0] _io_ca_T_1 = io_in_0 & io_in_2; // @[Compressor32.scala 22:25]
  wire [64:0] _io_ca_T_2 = _io_ca_T | _io_ca_T_1; // @[Compressor32.scala 22:20]
  wire [64:0] _io_ca_T_3 = io_in_1 & io_in_2; // @[Compressor32.scala 22:37]
  assign io_s = _io_s_T ^ io_in_2; // @[Compressor32.scala 21:17]
  assign io_ca = _io_ca_T_2 | _io_ca_T_3; // @[Compressor32.scala 22:32]
endmodule
module Multiplier19(
  input          clk_in1_p,
  input          clk_in1_n,
  input          reset,
  input          io_down_0,
  input          io_down_1,
  input  [64:0]  io_multiplicand,
  input  [64:0]  io_multiplier,
  input  [64:0]  io_addend,
  input          io_sub_vld,
  output [129:0] io_product
);
  clk_wiz_0 clk_wiz
   (
    // Clock out ports
    .clk_out1(clock),     		// output clk_out1
    // Clock in ports
    .clk_in1_p(clk_in1_p),    	// input clk_in1_p
    .clk_in1_n(clk_in1_n));    	// input clk_in1_n

`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [95:0] _RAND_14;
  reg [95:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire [64:0] boothCodeOutput_boothCodeUnit_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_1_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_1_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_2_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_2_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_3_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_3_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_4_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_4_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_5_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_5_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_6_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_6_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_7_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_7_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_8_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_8_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_9_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_9_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_10_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_10_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_11_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_11_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_12_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_12_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_13_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_13_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_14_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_14_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_15_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_15_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_16_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_16_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_17_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_17_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_18_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_18_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_19_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_19_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_20_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_20_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_21_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_21_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_22_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_22_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_23_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_23_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_24_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_24_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_25_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_25_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_26_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_26_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_27_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_27_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_28_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_28_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_29_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_29_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_30_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_30_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_31_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_31_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [64:0] boothCodeOutput_boothCodeUnit_32_io_A; // @[BoothCode.scala 66:31]
  wire [2:0] boothCodeOutput_boothCodeUnit_32_io_code; // @[BoothCode.scala 66:31]
  wire [65:0] boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_product; // @[BoothCode.scala 66:31]
  wire [1:0] boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_h; // @[BoothCode.scala 66:31]
  wire  boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_sn; // @[BoothCode.scala 66:31]
  wire [72:0] compressorOutLast_outs_compressor32_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_1_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_1_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_1_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_1_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_1_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_2_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_2_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_2_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_2_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_2_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_3_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_3_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_3_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_3_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_3_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_4_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_4_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_4_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_4_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_4_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_5_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_5_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_5_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_5_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_5_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_6_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_6_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_6_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_6_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_6_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_7_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_7_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_7_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_7_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_7_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_8_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_8_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_8_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_8_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_8_io_ca; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_9_io_in_0; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_9_io_in_1; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_9_io_in_2; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_9_io_s; // @[Compressor32.scala 42:44]
  wire [72:0] compressorOutLast_outs_compressor32_9_io_ca; // @[Compressor32.scala 42:44]
  wire [68:0] compressorOutLast_outs_compressor32_10_io_in_0; // @[Compressor32.scala 42:44]
  wire [68:0] compressorOutLast_outs_compressor32_10_io_in_1; // @[Compressor32.scala 42:44]
  wire [68:0] compressorOutLast_outs_compressor32_10_io_in_2; // @[Compressor32.scala 42:44]
  wire [68:0] compressorOutLast_outs_compressor32_10_io_s; // @[Compressor32.scala 42:44]
  wire [68:0] compressorOutLast_outs_compressor32_10_io_ca; // @[Compressor32.scala 42:44]
  wire [74:0] compressorOutLast_outs_compressor42_io_p_0; // @[Compressor42.scala 50:44]
  wire [74:0] compressorOutLast_outs_compressor42_io_p_1; // @[Compressor42.scala 50:44]
  wire [74:0] compressorOutLast_outs_compressor42_io_p_2; // @[Compressor42.scala 50:44]
  wire [74:0] compressorOutLast_outs_compressor42_io_p_3; // @[Compressor42.scala 50:44]
  wire [74:0] compressorOutLast_outs_compressor42_io_s; // @[Compressor42.scala 50:44]
  wire [74:0] compressorOutLast_outs_compressor42_io_ca; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_1_io_p_0; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_1_io_p_1; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_1_io_p_2; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_1_io_p_3; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_1_io_s; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_1_io_ca; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_2_io_p_0; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_2_io_p_1; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_2_io_p_2; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_2_io_p_3; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_2_io_s; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_2_io_ca; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_3_io_p_0; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_3_io_p_1; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_3_io_p_2; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_3_io_p_3; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_3_io_s; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_3_io_ca; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_4_io_p_0; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_4_io_p_1; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_4_io_p_2; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_4_io_p_3; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_4_io_s; // @[Compressor42.scala 50:44]
  wire [79:0] compressorOutLast_outs_compressor42_4_io_ca; // @[Compressor42.scala 50:44]
  wire [75:0] compressorOutLast_outs_compressor42_5_io_p_0; // @[Compressor42.scala 50:44]
  wire [75:0] compressorOutLast_outs_compressor42_5_io_p_1; // @[Compressor42.scala 50:44]
  wire [75:0] compressorOutLast_outs_compressor42_5_io_p_2; // @[Compressor42.scala 50:44]
  wire [75:0] compressorOutLast_outs_compressor42_5_io_p_3; // @[Compressor42.scala 50:44]
  wire [75:0] compressorOutLast_outs_compressor42_5_io_s; // @[Compressor42.scala 50:44]
  wire [75:0] compressorOutLast_outs_compressor42_5_io_ca; // @[Compressor42.scala 50:44]
  wire [86:0] compressorOutLast_outs_compressor32_11_io_in_0; // @[Compressor32.scala 42:44]
  wire [86:0] compressorOutLast_outs_compressor32_11_io_in_1; // @[Compressor32.scala 42:44]
  wire [86:0] compressorOutLast_outs_compressor32_11_io_in_2; // @[Compressor32.scala 42:44]
  wire [86:0] compressorOutLast_outs_compressor32_11_io_s; // @[Compressor32.scala 42:44]
  wire [86:0] compressorOutLast_outs_compressor32_11_io_ca; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_12_io_in_0; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_12_io_in_1; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_12_io_in_2; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_12_io_s; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_12_io_ca; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_13_io_in_0; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_13_io_in_1; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_13_io_in_2; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_13_io_s; // @[Compressor32.scala 42:44]
  wire [91:0] compressorOutLast_outs_compressor32_13_io_ca; // @[Compressor32.scala 42:44]
  wire [87:0] compressorOutLast_outs_compressor32_14_io_in_0; // @[Compressor32.scala 42:44]
  wire [87:0] compressorOutLast_outs_compressor32_14_io_in_1; // @[Compressor32.scala 42:44]
  wire [87:0] compressorOutLast_outs_compressor32_14_io_in_2; // @[Compressor32.scala 42:44]
  wire [87:0] compressorOutLast_outs_compressor32_14_io_s; // @[Compressor32.scala 42:44]
  wire [87:0] compressorOutLast_outs_compressor32_14_io_ca; // @[Compressor32.scala 42:44]
  wire [114:0] compressorOutLast_outs_compressor32_15_io_in_0; // @[Compressor32.scala 42:44]
  wire [114:0] compressorOutLast_outs_compressor32_15_io_in_1; // @[Compressor32.scala 42:44]
  wire [114:0] compressorOutLast_outs_compressor32_15_io_in_2; // @[Compressor32.scala 42:44]
  wire [114:0] compressorOutLast_outs_compressor32_15_io_s; // @[Compressor32.scala 42:44]
  wire [114:0] compressorOutLast_outs_compressor32_15_io_ca; // @[Compressor32.scala 42:44]
  wire [100:0] compressorOutLast_outs_compressor32_16_io_in_0; // @[Compressor32.scala 42:44]
  wire [100:0] compressorOutLast_outs_compressor32_16_io_in_1; // @[Compressor32.scala 42:44]
  wire [100:0] compressorOutLast_outs_compressor32_16_io_in_2; // @[Compressor32.scala 42:44]
  wire [100:0] compressorOutLast_outs_compressor32_16_io_s; // @[Compressor32.scala 42:44]
  wire [100:0] compressorOutLast_outs_compressor32_16_io_ca; // @[Compressor32.scala 42:44]
  wire [125:0] compressorOutLast_outs_compressor42_6_io_p_0; // @[Compressor42.scala 50:44]
  wire [125:0] compressorOutLast_outs_compressor42_6_io_p_1; // @[Compressor42.scala 50:44]
  wire [125:0] compressorOutLast_outs_compressor42_6_io_p_2; // @[Compressor42.scala 50:44]
  wire [125:0] compressorOutLast_outs_compressor42_6_io_p_3; // @[Compressor42.scala 50:44]
  wire [125:0] compressorOutLast_outs_compressor42_6_io_s; // @[Compressor42.scala 50:44]
  wire [125:0] compressorOutLast_outs_compressor42_6_io_ca; // @[Compressor42.scala 50:44]
  wire [132:0] compressorOutLast_outs_compressor42_7_io_p_0; // @[Compressor42.scala 50:44]
  wire [132:0] compressorOutLast_outs_compressor42_7_io_p_1; // @[Compressor42.scala 50:44]
  wire [132:0] compressorOutLast_outs_compressor42_7_io_p_2; // @[Compressor42.scala 50:44]
  wire [132:0] compressorOutLast_outs_compressor42_7_io_p_3; // @[Compressor42.scala 50:44]
  wire [132:0] compressorOutLast_outs_compressor42_7_io_s; // @[Compressor42.scala 50:44]
  wire [132:0] compressorOutLast_outs_compressor42_7_io_ca; // @[Compressor42.scala 50:44]
  wire [64:0] compressor32Out_compressor32_io_in_0; // @[Compressor32.scala 42:44]
  wire [64:0] compressor32Out_compressor32_io_in_1; // @[Compressor32.scala 42:44]
  wire [64:0] compressor32Out_compressor32_io_in_2; // @[Compressor32.scala 42:44]
  wire [64:0] compressor32Out_compressor32_io_s; // @[Compressor32.scala 42:44]
  wire [64:0] compressor32Out_compressor32_io_ca; // @[Compressor32.scala 42:44]
  wire [64:0] _multiplicand_not_T_2 = ~io_multiplicand; // @[Multiplier.scala 23:44]
  wire [64:0] _boothCodeOutput_T = io_multiplier; // @[Multiplier.scala 29:92]
  wire [63:0] partProductLast = io_sub_vld ? io_multiplier[63:0] : 64'h0; // @[Multiplier.scala 34:20 35:21 37:21]
  wire  boothCodeOutput_0_sn = boothCodeOutput_boothCodeUnit_io_boothCodeOutput_sn; // @[BoothCode.scala 83:{14,14}]
  wire  _partProducts_pProduct_0_value_T = ~boothCodeOutput_0_sn; // @[BCOutput2PProduct.scala 14:58]
  wire [65:0] boothCodeOutput_0_product = boothCodeOutput_boothCodeUnit_io_boothCodeOutput_product; // @[BoothCode.scala 83:{14,14}]
  wire [66:0] partProducts_pProduct_0_value_lo = {_partProducts_pProduct_0_value_T,boothCodeOutput_0_product}; // @[Cat.scala 31:58]
  wire [1:0] partProducts_pProduct_0_value_hi = {boothCodeOutput_0_sn,_partProducts_pProduct_0_value_T}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_1_sn = boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_1_product = boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [66:0] partProducts_pProduct_1_value_hi = {boothCodeOutput_1_sn,boothCodeOutput_1_product}; // @[Cat.scala 31:58]
  wire [1:0] boothCodeOutput_0_h = boothCodeOutput_boothCodeUnit_io_boothCodeOutput_h; // @[BoothCode.scala 83:{14,14}]
  wire  boothCodeOutput_2_sn = boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_2_product = boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_1_h = boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_2_value = {boothCodeOutput_2_sn,boothCodeOutput_2_product,boothCodeOutput_1_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_3_sn = boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_3_product = boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_2_h = boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_4_sn = boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_4_product = boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_3_h = boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_4_value = {boothCodeOutput_4_sn,boothCodeOutput_4_product,boothCodeOutput_3_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_5_sn = boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_5_product = boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_4_h = boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_5_value = {boothCodeOutput_5_sn,boothCodeOutput_5_product,boothCodeOutput_4_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_6_sn = boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_6_product = boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_5_h = boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_7_sn = boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_7_product = boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_6_h = boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_7_value = {boothCodeOutput_7_sn,boothCodeOutput_7_product,boothCodeOutput_6_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_8_sn = boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_8_product = boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_7_h = boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_8_value = {boothCodeOutput_8_sn,boothCodeOutput_8_product,boothCodeOutput_7_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_9_sn = boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_9_product = boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_8_h = boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_10_sn = boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_10_product = boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_9_h = boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_10_value = {boothCodeOutput_10_sn,boothCodeOutput_10_product,boothCodeOutput_9_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_11_sn = boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_11_product = boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_10_h = boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_11_value = {boothCodeOutput_11_sn,boothCodeOutput_11_product,boothCodeOutput_10_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_12_sn = boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_12_product = boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_11_h = boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_13_sn = boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_13_product = boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_12_h = boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_13_value = {boothCodeOutput_13_sn,boothCodeOutput_13_product,boothCodeOutput_12_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_14_sn = boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_14_product = boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_13_h = boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_14_value = {boothCodeOutput_14_sn,boothCodeOutput_14_product,boothCodeOutput_13_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_15_sn = boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_15_product = boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_14_h = boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_16_sn = boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_16_product = boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_15_h = boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_16_value = {boothCodeOutput_16_sn,boothCodeOutput_16_product,boothCodeOutput_15_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_17_sn = boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_17_product = boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_16_h = boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_17_value = {boothCodeOutput_17_sn,boothCodeOutput_17_product,boothCodeOutput_16_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_18_sn = boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_18_product = boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_17_h = boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_19_sn = boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_19_product = boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_18_h = boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_19_value = {boothCodeOutput_19_sn,boothCodeOutput_19_product,boothCodeOutput_18_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_20_sn = boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_20_product = boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_19_h = boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_20_value = {boothCodeOutput_20_sn,boothCodeOutput_20_product,boothCodeOutput_19_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_21_sn = boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_21_product = boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_20_h = boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_22_sn = boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_22_product = boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_21_h = boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_22_value = {boothCodeOutput_22_sn,boothCodeOutput_22_product,boothCodeOutput_21_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_23_sn = boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_23_product = boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_22_h = boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_23_value = {boothCodeOutput_23_sn,boothCodeOutput_23_product,boothCodeOutput_22_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_24_sn = boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_24_product = boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_23_h = boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_25_sn = boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_25_product = boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_24_h = boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_25_value = {boothCodeOutput_25_sn,boothCodeOutput_25_product,boothCodeOutput_24_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_26_sn = boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_26_product = boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_25_h = boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_26_value = {boothCodeOutput_26_sn,boothCodeOutput_26_product,boothCodeOutput_25_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_27_sn = boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_27_product = boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_26_h = boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_28_sn = boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_28_product = boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_27_h = boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_28_value = {boothCodeOutput_28_sn,boothCodeOutput_28_product,boothCodeOutput_27_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_29_sn = boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_29_product = boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_28_h = boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_29_value = {boothCodeOutput_29_sn,boothCodeOutput_29_product,boothCodeOutput_28_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_30_sn = boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_30_product = boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_29_h = boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire  boothCodeOutput_31_sn = boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_sn; // @[BoothCode.scala 87:{14,14}]
  wire [65:0] boothCodeOutput_31_product = boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_product; // @[BoothCode.scala 87:{14,14}]
  wire [1:0] boothCodeOutput_30_h = boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] partProducts_pProduct_31_value = {boothCodeOutput_31_sn,boothCodeOutput_31_product,boothCodeOutput_30_h}; // @[Cat.scala 31:58]
  wire  boothCodeOutput_32_sn = boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_sn; // @[BoothCode.scala 91:{14,14}]
  wire [65:0] boothCodeOutput_32_product = boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_product; // @[BoothCode.scala 91:{14,14}]
  wire [1:0] boothCodeOutput_31_h = boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_h; // @[BoothCode.scala 87:{14,14}]
  wire [68:0] _partProducts_valueLen_value_T = {boothCodeOutput_32_sn,boothCodeOutput_32_product,boothCodeOutput_31_h}; // @[Cat.scala 31:58]
  wire [1:0] boothCodeOutput_32_h = boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_h; // @[BoothCode.scala 91:{14,14}]
  wire  _partProducts_valueLenPlus2_value_T_1 = ~partProductLast[63]; // @[BCOutput2PProduct.scala 35:81]
  wire [65:0] partProducts_34_value = {_partProducts_valueLenPlus2_value_T_1,partProductLast[63],partProductLast}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_1 = {boothCodeOutput_30_sn,boothCodeOutput_30_product,
    boothCodeOutput_29_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_3 = {boothCodeOutput_27_sn,boothCodeOutput_27_product,
    boothCodeOutput_26_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_5 = {boothCodeOutput_24_sn,boothCodeOutput_24_product,
    boothCodeOutput_23_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_7 = {boothCodeOutput_21_sn,boothCodeOutput_21_product,
    boothCodeOutput_20_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_9 = {boothCodeOutput_18_sn,boothCodeOutput_18_product,
    boothCodeOutput_17_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_11 = {boothCodeOutput_15_sn,boothCodeOutput_15_product,
    boothCodeOutput_14_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_13 = {boothCodeOutput_12_sn,boothCodeOutput_12_product,
    boothCodeOutput_11_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_15 = {boothCodeOutput_9_sn,boothCodeOutput_9_product,
    boothCodeOutput_8_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_17 = {boothCodeOutput_6_sn,boothCodeOutput_6_product,
    boothCodeOutput_5_h,2'h0}; // @[Cat.scala 31:58]
  wire [70:0] _compressorOutLast_outs_compressor32_io_in_1_T_19 = {boothCodeOutput_3_sn,boothCodeOutput_3_product,
    boothCodeOutput_2_h,2'h0}; // @[Cat.scala 31:58]
  wire [67:0] partProducts_32_value = _partProducts_valueLen_value_T[67:0]; // @[BCOutput2PProduct.scala 25:24 26:20]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_1_T_1 = {partProducts_32_value,6'h0}; // @[Cat.scala 31:58]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_2_T_1 = {61'h1555555555555554,4'hf,boothCodeOutput_32_h[0],8'h0}
    ; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_ca_value = compressorOutLast_outs_compressor32_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_3_T = {compressorOutLast_outs_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_2_ca_value = compressorOutLast_outs_compressor32_2_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_1_T_2 = {compressorOutLast_outs_2_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_1_s_value = compressorOutLast_outs_compressor32_1_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [78:0] _compressorOutLast_outs_compressor42_io_p_2_T_3 = {compressorOutLast_outs_1_s_value,6'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_1_ca_value = compressorOutLast_outs_compressor32_1_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [72:0] compressorOutLast_outs_4_ca_value = compressorOutLast_outs_compressor32_4_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_1_T_3 = {compressorOutLast_outs_4_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_3_s_value = compressorOutLast_outs_compressor32_3_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [78:0] _compressorOutLast_outs_compressor42_io_p_2_T_5 = {compressorOutLast_outs_3_s_value,6'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_3_ca_value = compressorOutLast_outs_compressor32_3_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [72:0] compressorOutLast_outs_6_ca_value = compressorOutLast_outs_compressor32_6_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_1_T_4 = {compressorOutLast_outs_6_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_5_s_value = compressorOutLast_outs_compressor32_5_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [78:0] _compressorOutLast_outs_compressor42_io_p_2_T_7 = {compressorOutLast_outs_5_s_value,6'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_5_ca_value = compressorOutLast_outs_compressor32_5_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [72:0] compressorOutLast_outs_8_ca_value = compressorOutLast_outs_compressor32_8_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [73:0] _compressorOutLast_outs_compressor42_io_p_1_T_5 = {compressorOutLast_outs_8_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_7_s_value = compressorOutLast_outs_compressor32_7_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [78:0] _compressorOutLast_outs_compressor42_io_p_2_T_9 = {compressorOutLast_outs_7_s_value,6'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_7_ca_value = compressorOutLast_outs_compressor32_7_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [68:0] compressorOutLast_outs_10_ca_value = compressorOutLast_outs_compressor32_10_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [69:0] _compressorOutLast_outs_compressor42_io_p_1_T_6 = {compressorOutLast_outs_10_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_9_s_value = compressorOutLast_outs_compressor32_9_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [74:0] _compressorOutLast_outs_compressor42_io_p_2_T_11 = {compressorOutLast_outs_9_s_value,2'h0}; // @[Cat.scala 31:58]
  wire [72:0] compressorOutLast_outs_9_ca_value = compressorOutLast_outs_compressor32_9_io_ca; // @[Compressor32.scala 49:50 51:31]
  reg [75:0] compressorOutLast_regC; // @[Compressor.scala 109:29]
  wire [75:0] compressorOutLast_outs_16_s_value = compressorOutLast_outs_compressor42_5_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [75:0] compressorOutLast_regC_1; // @[Compressor.scala 109:29]
  wire [75:0] compressorOutLast_outs_16_ca_value = compressorOutLast_outs_compressor42_5_io_ca; // @[Compressor42.scala 57:50 59:31]
  reg [79:0] compressorOutLast_regC_2; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_15_s_value = compressorOutLast_outs_compressor42_4_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [79:0] compressorOutLast_regC_3; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_15_ca_value = compressorOutLast_outs_compressor42_4_io_ca; // @[Compressor42.scala 57:50 59:31]
  reg [79:0] compressorOutLast_regC_4; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_14_s_value = compressorOutLast_outs_compressor42_3_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [79:0] compressorOutLast_regC_5; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_14_ca_value = compressorOutLast_outs_compressor42_3_io_ca; // @[Compressor42.scala 57:50 59:31]
  reg [79:0] compressorOutLast_regC_6; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_13_s_value = compressorOutLast_outs_compressor42_2_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [79:0] compressorOutLast_regC_7; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_13_ca_value = compressorOutLast_outs_compressor42_2_io_ca; // @[Compressor42.scala 57:50 59:31]
  reg [79:0] compressorOutLast_regC_8; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_12_s_value = compressorOutLast_outs_compressor42_1_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [79:0] compressorOutLast_regC_9; // @[Compressor.scala 109:29]
  wire [79:0] compressorOutLast_outs_12_ca_value = compressorOutLast_outs_compressor42_1_io_ca; // @[Compressor42.scala 57:50 59:31]
  reg [74:0] compressorOutLast_regC_10; // @[Compressor.scala 109:29]
  wire [74:0] compressorOutLast_outs_11_s_value = compressorOutLast_outs_compressor42_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [74:0] compressorOutLast_regC_11; // @[Compressor.scala 109:29]
  wire [74:0] compressorOutLast_outs_11_ca_value = compressorOutLast_outs_compressor42_io_ca; // @[Compressor42.scala 57:50 59:31]
  wire [85:0] _compressorOutLast_outs_compressor32_io_in_1_T_21 = {compressorOutLast_regC_10,11'h0}; // @[Cat.scala 31:58]
  wire [80:0] _compressorOutLast_outs_compressor32_io_in_1_T_22 = {compressorOutLast_regC_7,1'h0}; // @[Cat.scala 31:58]
  wire [90:0] _compressorOutLast_outs_compressor32_io_in_1_T_24 = {compressorOutLast_regC_4,11'h0}; // @[Cat.scala 31:58]
  wire [76:0] _compressorOutLast_outs_compressor32_io_in_1_T_25 = {compressorOutLast_regC_1,1'h0}; // @[Cat.scala 31:58]
  wire [91:0] compressorOutLast_outs_18_s_value = compressorOutLast_outs_compressor32_12_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [113:0] _compressorOutLast_outs_compressor32_io_in_1_T_27 = {compressorOutLast_outs_18_s_value,22'h0}; // @[Cat.scala 31:58]
  wire [91:0] compressorOutLast_outs_18_ca_value = compressorOutLast_outs_compressor32_12_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [87:0] compressorOutLast_outs_20_ca_value = compressorOutLast_outs_compressor32_14_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [88:0] _compressorOutLast_outs_compressor32_io_in_1_T_28 = {compressorOutLast_outs_20_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [91:0] compressorOutLast_outs_19_s_value = compressorOutLast_outs_compressor32_13_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [100:0] compressorOutLast_outs_22_ca_value = compressorOutLast_outs_compressor32_16_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [101:0] _compressorOutLast_outs_compressor42_io_p_1_T_7 = {compressorOutLast_outs_22_ca_value,1'h0}; // @[Cat.scala 31:58]
  wire [114:0] compressorOutLast_outs_21_s_value = compressorOutLast_outs_compressor32_15_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [124:0] _compressorOutLast_outs_compressor42_io_p_2_T_13 = {compressorOutLast_outs_21_s_value,10'h0}; // @[Cat.scala 31:58]
  wire [114:0] compressorOutLast_outs_21_ca_value = compressorOutLast_outs_compressor32_15_io_ca; // @[Compressor32.scala 49:50 51:31]
  reg [125:0] compressorOutLast_regC_12; // @[Compressor.scala 109:29]
  wire [125:0] compressorOutLast_outs_23_s_value = compressorOutLast_outs_compressor42_6_io_s; // @[Compressor42.scala 57:50 58:30]
  reg [125:0] compressorOutLast_regC_13; // @[Compressor.scala 109:29]
  wire [125:0] compressorOutLast_outs_23_ca_value = compressorOutLast_outs_compressor42_6_io_ca; // @[Compressor42.scala 57:50 59:31]
  reg [86:0] compressorOutLast_regC_14; // @[Compressor.scala 109:29]
  wire [86:0] compressorOutLast_outs_17_s_value = compressorOutLast_outs_compressor32_11_io_s; // @[Compressor32.scala 49:50 50:30]
  reg [86:0] compressorOutLast_regC_15; // @[Compressor.scala 109:29]
  wire [86:0] compressorOutLast_outs_17_ca_value = compressorOutLast_outs_compressor32_11_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [126:0] _compressorOutLast_outs_compressor42_io_p_1_T_8 = {compressorOutLast_regC_13,1'h0}; // @[Cat.scala 31:58]
  wire [131:0] _compressorOutLast_outs_compressor42_io_p_2_T_15 = {compressorOutLast_regC_14,45'h0}; // @[Cat.scala 31:58]
  wire [132:0] compressorOutLast_outs_24_s_value = compressorOutLast_outs_compressor42_7_io_s; // @[Compressor42.scala 57:50 58:30]
  wire [129:0] sum = compressorOutLast_outs_24_s_value[129:0]; // @[Multiplier.scala 55:23 58:7]
  wire [63:0] compressor32Out_compressor32In_0_value = sum[63:0]; // @[AddAddend.scala 8:35]
  wire [132:0] compressorOutLast_outs_24_ca_value = compressorOutLast_outs_compressor42_7_io_ca; // @[Compressor42.scala 57:50 59:31]
  wire [129:0] carry = compressorOutLast_outs_24_ca_value[129:0]; // @[Multiplier.scala 56:25 59:9]
  wire [63:0] compressor32Out_compressor32In_1_value = carry[63:0]; // @[AddAddend.scala 10:37]
  wire [63:0] compressor32Out_compressor32In_2_value = io_addend[63:0]; // @[AddAddend.scala 12:39]
  wire [130:0] _productMult_T = {carry, 1'h0}; // @[Multiplier.scala 71:25]
  wire [130:0] _GEN_19 = {{1'd0}, sum}; // @[Multiplier.scala 71:38]
  wire [130:0] _productMult_T_2 = _productMult_T + _GEN_19; // @[Multiplier.scala 71:38]
  wire [64:0] compressor32Out_ca_value = compressor32Out_compressor32_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [65:0] _productMultAdd_T = {compressor32Out_ca_value, 1'h0}; // @[Multiplier.scala 72:47]
  wire [64:0] compressor32Out_s_value = compressor32Out_compressor32_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [65:0] _GEN_20 = {{1'd0}, compressor32Out_s_value}; // @[Multiplier.scala 72:60]
  wire [65:0] _productMultAdd_T_2 = _productMultAdd_T + _GEN_20; // @[Multiplier.scala 72:60]
  wire [129:0] productMult = _productMult_T_2[129:0]; // @[Multiplier.scala 69:31 71:15]
  wire [63:0] productMultAdd = _productMultAdd_T_2[63:0]; // @[Multiplier.scala 70:34 72:18]
  wire [72:0] compressorOutLast_outs_s_value = compressorOutLast_outs_compressor32_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [72:0] compressorOutLast_outs_2_s_value = compressorOutLast_outs_compressor32_2_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [72:0] compressorOutLast_outs_4_s_value = compressorOutLast_outs_compressor32_4_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [72:0] compressorOutLast_outs_6_s_value = compressorOutLast_outs_compressor32_6_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [72:0] compressorOutLast_outs_8_s_value = compressorOutLast_outs_compressor32_8_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [68:0] compressorOutLast_outs_10_s_value = compressorOutLast_outs_compressor32_10_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [91:0] compressorOutLast_outs_19_ca_value = compressorOutLast_outs_compressor32_13_io_ca; // @[Compressor32.scala 49:50 51:31]
  wire [87:0] compressorOutLast_outs_20_s_value = compressorOutLast_outs_compressor32_14_io_s; // @[Compressor32.scala 49:50 50:30]
  wire [100:0] compressorOutLast_outs_22_s_value = compressorOutLast_outs_compressor32_16_io_s; // @[Compressor32.scala 49:50 50:30]
  BoothCodeUnit boothCodeOutput_boothCodeUnit ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_1 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_1_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_1_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_1_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_2 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_2_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_2_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_2_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_3 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_3_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_3_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_3_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_4 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_4_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_4_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_4_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_5 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_5_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_5_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_5_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_6 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_6_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_6_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_6_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_7 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_7_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_7_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_7_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_8 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_8_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_8_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_8_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_9 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_9_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_9_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_9_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_10 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_10_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_10_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_10_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_11 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_11_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_11_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_11_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_12 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_12_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_12_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_12_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_13 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_13_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_13_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_13_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_14 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_14_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_14_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_14_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_15 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_15_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_15_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_15_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_16 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_16_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_16_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_16_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_17 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_17_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_17_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_17_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_18 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_18_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_18_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_18_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_19 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_19_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_19_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_19_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_20 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_20_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_20_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_20_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_21 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_21_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_21_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_21_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_22 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_22_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_22_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_22_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_23 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_23_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_23_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_23_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_24 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_24_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_24_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_24_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_25 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_25_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_25_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_25_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_26 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_26_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_26_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_26_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_27 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_27_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_27_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_27_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_28 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_28_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_28_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_28_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_29 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_29_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_29_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_29_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_30 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_30_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_30_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_30_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_31 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_31_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_31_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_31_io_boothCodeOutput_sn)
  );
  BoothCodeUnit boothCodeOutput_boothCodeUnit_32 ( // @[BoothCode.scala 66:31]
    .io_A(boothCodeOutput_boothCodeUnit_32_io_A),
    .io_code(boothCodeOutput_boothCodeUnit_32_io_code),
    .io_boothCodeOutput_product(boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_product),
    .io_boothCodeOutput_h(boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_h),
    .io_boothCodeOutput_sn(boothCodeOutput_boothCodeUnit_32_io_boothCodeOutput_sn)
  );
  Compressor32 compressorOutLast_outs_compressor32 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_io_s),
    .io_ca(compressorOutLast_outs_compressor32_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_1 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_1_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_1_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_1_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_1_io_s),
    .io_ca(compressorOutLast_outs_compressor32_1_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_2 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_2_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_2_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_2_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_2_io_s),
    .io_ca(compressorOutLast_outs_compressor32_2_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_3 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_3_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_3_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_3_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_3_io_s),
    .io_ca(compressorOutLast_outs_compressor32_3_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_4 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_4_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_4_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_4_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_4_io_s),
    .io_ca(compressorOutLast_outs_compressor32_4_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_5 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_5_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_5_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_5_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_5_io_s),
    .io_ca(compressorOutLast_outs_compressor32_5_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_6 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_6_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_6_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_6_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_6_io_s),
    .io_ca(compressorOutLast_outs_compressor32_6_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_7 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_7_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_7_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_7_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_7_io_s),
    .io_ca(compressorOutLast_outs_compressor32_7_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_8 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_8_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_8_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_8_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_8_io_s),
    .io_ca(compressorOutLast_outs_compressor32_8_io_ca)
  );
  Compressor32 compressorOutLast_outs_compressor32_9 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_9_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_9_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_9_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_9_io_s),
    .io_ca(compressorOutLast_outs_compressor32_9_io_ca)
  );
  Compressor32_10 compressorOutLast_outs_compressor32_10 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_10_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_10_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_10_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_10_io_s),
    .io_ca(compressorOutLast_outs_compressor32_10_io_ca)
  );
  Compressor42 compressorOutLast_outs_compressor42 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_io_s),
    .io_ca(compressorOutLast_outs_compressor42_io_ca)
  );
  Compressor42_1 compressorOutLast_outs_compressor42_1 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_1_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_1_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_1_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_1_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_1_io_s),
    .io_ca(compressorOutLast_outs_compressor42_1_io_ca)
  );
  Compressor42_1 compressorOutLast_outs_compressor42_2 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_2_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_2_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_2_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_2_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_2_io_s),
    .io_ca(compressorOutLast_outs_compressor42_2_io_ca)
  );
  Compressor42_1 compressorOutLast_outs_compressor42_3 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_3_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_3_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_3_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_3_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_3_io_s),
    .io_ca(compressorOutLast_outs_compressor42_3_io_ca)
  );
  Compressor42_1 compressorOutLast_outs_compressor42_4 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_4_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_4_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_4_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_4_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_4_io_s),
    .io_ca(compressorOutLast_outs_compressor42_4_io_ca)
  );
  Compressor42_5 compressorOutLast_outs_compressor42_5 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_5_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_5_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_5_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_5_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_5_io_s),
    .io_ca(compressorOutLast_outs_compressor42_5_io_ca)
  );
  Compressor32_11 compressorOutLast_outs_compressor32_11 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_11_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_11_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_11_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_11_io_s),
    .io_ca(compressorOutLast_outs_compressor32_11_io_ca)
  );
  Compressor32_12 compressorOutLast_outs_compressor32_12 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_12_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_12_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_12_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_12_io_s),
    .io_ca(compressorOutLast_outs_compressor32_12_io_ca)
  );
  Compressor32_12 compressorOutLast_outs_compressor32_13 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_13_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_13_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_13_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_13_io_s),
    .io_ca(compressorOutLast_outs_compressor32_13_io_ca)
  );
  Compressor32_14 compressorOutLast_outs_compressor32_14 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_14_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_14_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_14_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_14_io_s),
    .io_ca(compressorOutLast_outs_compressor32_14_io_ca)
  );
  Compressor32_15 compressorOutLast_outs_compressor32_15 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_15_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_15_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_15_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_15_io_s),
    .io_ca(compressorOutLast_outs_compressor32_15_io_ca)
  );
  Compressor32_16 compressorOutLast_outs_compressor32_16 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressorOutLast_outs_compressor32_16_io_in_0),
    .io_in_1(compressorOutLast_outs_compressor32_16_io_in_1),
    .io_in_2(compressorOutLast_outs_compressor32_16_io_in_2),
    .io_s(compressorOutLast_outs_compressor32_16_io_s),
    .io_ca(compressorOutLast_outs_compressor32_16_io_ca)
  );
  Compressor42_6 compressorOutLast_outs_compressor42_6 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_6_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_6_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_6_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_6_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_6_io_s),
    .io_ca(compressorOutLast_outs_compressor42_6_io_ca)
  );
  Compressor42_7 compressorOutLast_outs_compressor42_7 ( // @[Compressor42.scala 50:44]
    .io_p_0(compressorOutLast_outs_compressor42_7_io_p_0),
    .io_p_1(compressorOutLast_outs_compressor42_7_io_p_1),
    .io_p_2(compressorOutLast_outs_compressor42_7_io_p_2),
    .io_p_3(compressorOutLast_outs_compressor42_7_io_p_3),
    .io_s(compressorOutLast_outs_compressor42_7_io_s),
    .io_ca(compressorOutLast_outs_compressor42_7_io_ca)
  );
  Compressor32_17 compressor32Out_compressor32 ( // @[Compressor32.scala 42:44]
    .io_in_0(compressor32Out_compressor32_io_in_0),
    .io_in_1(compressor32Out_compressor32_io_in_1),
    .io_in_2(compressor32Out_compressor32_io_in_2),
    .io_s(compressor32Out_compressor32_io_s),
    .io_ca(compressor32Out_compressor32_io_ca)
  );
  assign io_product = {productMult[129:64],productMultAdd}; // @[Multiplier.scala 74:67]
  assign boothCodeOutput_boothCodeUnit_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_io_code = {_boothCodeOutput_T[1:0],1'h0}; // @[Cat.scala 31:58]
  assign boothCodeOutput_boothCodeUnit_1_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_1_io_code = _boothCodeOutput_T[3:1]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_2_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_2_io_code = _boothCodeOutput_T[5:3]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_3_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_3_io_code = _boothCodeOutput_T[7:5]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_4_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_4_io_code = _boothCodeOutput_T[9:7]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_5_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_5_io_code = _boothCodeOutput_T[11:9]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_6_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_6_io_code = _boothCodeOutput_T[13:11]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_7_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_7_io_code = _boothCodeOutput_T[15:13]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_8_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_8_io_code = _boothCodeOutput_T[17:15]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_9_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_9_io_code = _boothCodeOutput_T[19:17]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_10_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_10_io_code = _boothCodeOutput_T[21:19]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_11_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_11_io_code = _boothCodeOutput_T[23:21]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_12_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_12_io_code = _boothCodeOutput_T[25:23]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_13_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_13_io_code = _boothCodeOutput_T[27:25]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_14_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_14_io_code = _boothCodeOutput_T[29:27]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_15_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_15_io_code = _boothCodeOutput_T[31:29]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_16_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_16_io_code = _boothCodeOutput_T[33:31]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_17_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_17_io_code = _boothCodeOutput_T[35:33]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_18_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_18_io_code = _boothCodeOutput_T[37:35]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_19_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_19_io_code = _boothCodeOutput_T[39:37]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_20_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_20_io_code = _boothCodeOutput_T[41:39]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_21_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_21_io_code = _boothCodeOutput_T[43:41]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_22_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_22_io_code = _boothCodeOutput_T[45:43]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_23_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_23_io_code = _boothCodeOutput_T[47:45]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_24_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_24_io_code = _boothCodeOutput_T[49:47]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_25_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_25_io_code = _boothCodeOutput_T[51:49]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_26_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_26_io_code = _boothCodeOutput_T[53:51]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_27_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_27_io_code = _boothCodeOutput_T[55:53]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_28_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_28_io_code = _boothCodeOutput_T[57:55]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_29_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_29_io_code = _boothCodeOutput_T[59:57]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_30_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_30_io_code = _boothCodeOutput_T[61:59]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_31_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_31_io_code = _boothCodeOutput_T[63:61]; // @[BoothCode.scala 87:78]
  assign boothCodeOutput_boothCodeUnit_32_io_A = io_sub_vld ? _multiplicand_not_T_2 : io_multiplicand; // @[Multiplier.scala 22:20 23:22 25:22]
  assign boothCodeOutput_boothCodeUnit_32_io_code = {_boothCodeOutput_T[64],_boothCodeOutput_T[64:63]}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_io_in_0 = {{4'd0}, partProducts_pProduct_29_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_1}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_io_in_2 = {partProducts_pProduct_31_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_1_io_in_0 = {{4'd0}, partProducts_pProduct_26_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_1_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_3}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_1_io_in_2 = {partProducts_pProduct_28_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_2_io_in_0 = {{4'd0}, partProducts_pProduct_23_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_2_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_5}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_2_io_in_2 = {partProducts_pProduct_25_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_3_io_in_0 = {{4'd0}, partProducts_pProduct_20_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_3_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_7}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_3_io_in_2 = {partProducts_pProduct_22_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_4_io_in_0 = {{4'd0}, partProducts_pProduct_17_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_4_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_9}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_4_io_in_2 = {partProducts_pProduct_19_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_5_io_in_0 = {{4'd0}, partProducts_pProduct_14_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_5_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_11}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_5_io_in_2 = {partProducts_pProduct_16_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_6_io_in_0 = {{4'd0}, partProducts_pProduct_11_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_6_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_13}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_6_io_in_2 = {partProducts_pProduct_13_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_7_io_in_0 = {{4'd0}, partProducts_pProduct_8_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_7_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_15}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_7_io_in_2 = {partProducts_pProduct_10_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_8_io_in_0 = {{4'd0}, partProducts_pProduct_5_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_8_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_17}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_8_io_in_2 = {partProducts_pProduct_7_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_9_io_in_0 = {{4'd0}, partProducts_pProduct_2_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_9_io_in_1 = {{2'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_19}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_9_io_in_2 = {partProducts_pProduct_4_value,4'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_10_io_in_0 = {{3'd0}, partProducts_34_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_10_io_in_1 = {partProducts_pProduct_0_value_hi,
    partProducts_pProduct_0_value_lo}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_10_io_in_2 = {partProducts_pProduct_1_value_hi,boothCodeOutput_0_h}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_io_p_0 = {{2'd0}, compressorOutLast_outs_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_io_p_1 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_1}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_1}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_io_p_3 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_3_T}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_1_io_p_0 = {{7'd0}, compressorOutLast_outs_2_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_1_io_p_1 = {{6'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_2}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_1_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_3}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_1_io_p_3 = {compressorOutLast_outs_1_ca_value,7'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_2_io_p_0 = {{7'd0}, compressorOutLast_outs_4_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_2_io_p_1 = {{6'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_3}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_2_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_5}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_2_io_p_3 = {compressorOutLast_outs_3_ca_value,7'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_3_io_p_0 = {{7'd0}, compressorOutLast_outs_6_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_3_io_p_1 = {{6'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_4}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_3_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_7}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_3_io_p_3 = {compressorOutLast_outs_5_ca_value,7'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_4_io_p_0 = {{7'd0}, compressorOutLast_outs_8_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_4_io_p_1 = {{6'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_5}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_4_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_9}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_4_io_p_3 = {compressorOutLast_outs_7_ca_value,7'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_5_io_p_0 = {{7'd0}, compressorOutLast_outs_10_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_5_io_p_1 = {{6'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_6}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_5_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_11}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_5_io_p_3 = {compressorOutLast_outs_9_ca_value,3'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_11_io_in_0 = {{7'd0}, compressorOutLast_regC_9}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_11_io_in_1 = {{1'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_21}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_11_io_in_2 = {compressorOutLast_regC_11,12'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_12_io_in_0 = {{12'd0}, compressorOutLast_regC_6}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_12_io_in_1 = {{11'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_22}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_12_io_in_2 = {compressorOutLast_regC_8,12'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_13_io_in_0 = {{12'd0}, compressorOutLast_regC_3}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_13_io_in_1 = {{1'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_24}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_13_io_in_2 = {compressorOutLast_regC_5,12'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_14_io_in_0 = {{12'd0}, compressorOutLast_regC}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_14_io_in_1 = {{11'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_25}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_14_io_in_2 = {compressorOutLast_regC_2,8'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_15_io_in_0 = {{23'd0}, compressorOutLast_outs_19_ca_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_15_io_in_1 = {{1'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_27}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_15_io_in_2 = {compressorOutLast_outs_18_ca_value,23'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor32_16_io_in_0 = {{13'd0}, compressorOutLast_outs_20_s_value}; // @[Compressor32.scala 45:51]
  assign compressorOutLast_outs_compressor32_16_io_in_1 = {{12'd0}, _compressorOutLast_outs_compressor32_io_in_1_T_28}; // @[Compressor32.scala 46:34]
  assign compressorOutLast_outs_compressor32_16_io_in_2 = {compressorOutLast_outs_19_s_value,9'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_6_io_p_0 = {{25'd0}, compressorOutLast_outs_22_s_value}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_6_io_p_1 = {{24'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_7}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_6_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_13}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_6_io_p_3 = {compressorOutLast_outs_21_ca_value,11'h0}; // @[Cat.scala 31:58]
  assign compressorOutLast_outs_compressor42_7_io_p_0 = {{7'd0}, compressorOutLast_regC_12}; // @[Compressor42.scala 53:50]
  assign compressorOutLast_outs_compressor42_7_io_p_1 = {{6'd0}, _compressorOutLast_outs_compressor42_io_p_1_T_8}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_7_io_p_2 = {{1'd0}, _compressorOutLast_outs_compressor42_io_p_2_T_15}; // @[Compressor42.scala 54:33]
  assign compressorOutLast_outs_compressor42_7_io_p_3 = {compressorOutLast_regC_15,46'h0}; // @[Cat.scala 31:58]
  assign compressor32Out_compressor32_io_in_0 = {{1'd0}, compressor32Out_compressor32In_0_value}; // @[Compressor32.scala 45:51]
  assign compressor32Out_compressor32_io_in_1 = {{1'd0}, compressor32Out_compressor32In_2_value}; // @[Compressor32.scala 45:51]
  assign compressor32Out_compressor32_io_in_2 = {compressor32Out_compressor32In_1_value,1'h0}; // @[Cat.scala 31:58]
  always @(posedge clock) begin
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC <= 76'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC <= compressorOutLast_outs_16_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_1 <= 76'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_1 <= compressorOutLast_outs_16_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_2 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_2 <= compressorOutLast_outs_15_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_3 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_3 <= compressorOutLast_outs_15_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_4 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_4 <= compressorOutLast_outs_14_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_5 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_5 <= compressorOutLast_outs_14_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_6 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_6 <= compressorOutLast_outs_13_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_7 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_7 <= compressorOutLast_outs_13_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_8 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_8 <= compressorOutLast_outs_12_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_9 <= 80'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_9 <= compressorOutLast_outs_12_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_10 <= 75'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_10 <= compressorOutLast_outs_11_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_11 <= 75'h0; // @[Compressor.scala 109:29]
    end else if (io_down_0) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_11 <= compressorOutLast_outs_11_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_12 <= 126'h0; // @[Compressor.scala 109:29]
    end else if (io_down_1) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_12 <= compressorOutLast_outs_23_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_13 <= 126'h0; // @[Compressor.scala 109:29]
    end else if (io_down_1) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_13 <= compressorOutLast_outs_23_ca_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_14 <= 87'h0; // @[Compressor.scala 109:29]
    end else if (io_down_1) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_14 <= compressorOutLast_outs_17_s_value; // @[Compressor.scala 112:18]
    end
    if (reset) begin // @[Compressor.scala 109:29]
      compressorOutLast_regC_15 <= 87'h0; // @[Compressor.scala 109:29]
    end else if (io_down_1) begin // @[Compressor.scala 111:28]
      compressorOutLast_regC_15 <= compressorOutLast_outs_17_ca_value; // @[Compressor.scala 112:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  compressorOutLast_regC = _RAND_0[75:0];
  _RAND_1 = {3{`RANDOM}};
  compressorOutLast_regC_1 = _RAND_1[75:0];
  _RAND_2 = {3{`RANDOM}};
  compressorOutLast_regC_2 = _RAND_2[79:0];
  _RAND_3 = {3{`RANDOM}};
  compressorOutLast_regC_3 = _RAND_3[79:0];
  _RAND_4 = {3{`RANDOM}};
  compressorOutLast_regC_4 = _RAND_4[79:0];
  _RAND_5 = {3{`RANDOM}};
  compressorOutLast_regC_5 = _RAND_5[79:0];
  _RAND_6 = {3{`RANDOM}};
  compressorOutLast_regC_6 = _RAND_6[79:0];
  _RAND_7 = {3{`RANDOM}};
  compressorOutLast_regC_7 = _RAND_7[79:0];
  _RAND_8 = {3{`RANDOM}};
  compressorOutLast_regC_8 = _RAND_8[79:0];
  _RAND_9 = {3{`RANDOM}};
  compressorOutLast_regC_9 = _RAND_9[79:0];
  _RAND_10 = {3{`RANDOM}};
  compressorOutLast_regC_10 = _RAND_10[74:0];
  _RAND_11 = {3{`RANDOM}};
  compressorOutLast_regC_11 = _RAND_11[74:0];
  _RAND_12 = {4{`RANDOM}};
  compressorOutLast_regC_12 = _RAND_12[125:0];
  _RAND_13 = {4{`RANDOM}};
  compressorOutLast_regC_13 = _RAND_13[125:0];
  _RAND_14 = {3{`RANDOM}};
  compressorOutLast_regC_14 = _RAND_14[86:0];
  _RAND_15 = {3{`RANDOM}};
  compressorOutLast_regC_15 = _RAND_15[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
